module  decimal_to_BCD_gold(D,Y);
input [9:0]D;
output [3:0]Y;
assign Y = (D==10'b0000000001)? 4'b0000 : 
(D== 10'b0000000010)?4'b0001:
(D==10'b0000000100)?4'b0010:
(D==10'b0000001000)?4'b0011:
(D==10'b0000010000)?4'b0100:
(D==10'b0000100000)?4'b0101:
(D==10'b0001000000)?4'b0110:
(D==10'b0010000000)?4'b0111:
(D==10'b0100000000)?4'b1000:
(D==10'b1000000000)?4'b1001:
4'b0000;
endmodule